module 
endmodule 
kncsin
skdnsd
