module 
endmodule 
kncsin
